library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

library work;
    use work.ethernet_frame_receiver_pkg.all;
    use work.ethernet_rx_ddio_pkg.all; 

package ethernet_frame_receiver_internal_pkg is

end package ethernet_frame_receiver_internal_pkg;


package body ethernet_frame_receiver_internal_pkg is


end package body ethernet_frame_receiver_internal_pkg;

