library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

-- entity network_protocol is
--     port (
--         network_protocol_clocks   : in network_protocol_clock_group;
--         network_protocol_data_in  : in network_protocol_data_input_group;
--         network_protocol_data_out : out network_protocol_data_output_group
--     );
-- end entity network_protocol;

architecture arch_internet_protocol of network_protocol is

    alias clock is network_protocol_clocks.clock;
    alias internet_protocol_data_in is network_protocol_data_in;
    alias internet_protocol_data_out is network_protocol_data_out;
    alias protocol_control is internet_protocol_data_in.protocol_control; 

    signal frame_ram_read_control_port : ram_read_control_group;
    signal shift_register : std_logic_vector(31 downto 0);
    signal ram_read_controller : ram_reader;
    signal ram_offset : natural range 0 to 2**11-1;
    signal header_offset : natural range 0 to 2**11-1;

------------------------------------------------------------------------ 
    signal udp_protocol_clocks   : network_protocol_clock_group;
    signal udp_protocol_data_in  : network_protocol_data_input_group;
    signal udp_protocol_data_out : network_protocol_data_output_group;
    signal udp_protocol_control  : protocol_control_record; 

begin

------------------------------------------------------------------------
    route_data_out : process(frame_ram_read_control_port, ram_offset, udp_protocol_data_out.frame_ram_read_control) 
    begin
        internet_protocol_data_out <= (
                                          frame_ram_read_control => frame_ram_read_control_port + udp_protocol_data_out.frame_ram_read_control,
                                          ram_offset => ram_offset
                                      );

    end process route_data_out;	
------------------------------------------------------------------------

    ip_header_processor : process(clock)
        
    begin
        if rising_edge(clock) then
            create_ram_read_controller(frame_ram_read_control_port, internet_protocol_data_in.frame_ram_output, ram_read_controller, shift_register); 
            init_protocol_control(udp_protocol_control);

            if protocol_control.protocol_processing_is_requested then
                load_ram_with_offset_to_shift_register(ram_controller                     => ram_read_controller,
                                                       start_address                      => protocol_control.protocol_start_address,
                                                       number_of_ram_addresses_to_be_read => 20);

                header_offset <= protocol_control.protocol_start_address;
            end if;

            if get_ram_address(internet_protocol_data_in.frame_ram_output) = header_offset+8 then
                if shift_register(7 downto 0) = x"11" then
                    ram_offset <= header_offset+8;
                    request_protocol_processing(udp_protocol_control, header_offset + 8);
                end if;
            end if;

        end if; --rising_edge
    end process ip_header_processor;	

------------------------------------------------------------------------ 
    udp_protocol_clocks <= (clock => clock);

    udp_protocol_data_in <= (frame_ram_output => internet_protocol_data_in.frame_ram_output, 
                                 protocol_control => udp_protocol_control);

    u_udp_protocol : entity work.network_protocol(arch_user_datagram_protocol)
    port map( udp_protocol_clocks  ,
              udp_protocol_data_in ,
              udp_protocol_data_out); 

------------------------------------------------------------------------ 
end arch_internet_protocol;
