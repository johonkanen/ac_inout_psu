library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

library math_library;
    use math_library.multiplier_pkg.all;
    use math_library.state_variable_pkg.all;
    use math_library.lcr_filter_model_pkg.all;

package inverter_model_pkg is

    type inverter_model_record is record
        inverter_multiplier : multiplier_record;
        inverter_lc_filter  : lcr_model_record;
        dc_link_voltage     : state_variable_record;

        duty_ratio                  : int18;
        dc_link_current             : int18;
        load_current                : int18;
        load_resistor_current       : int18;
        input_voltage               : int18;
        grid_inverter_state_counter : natural range 0 to 7;
    end record;

    constant init_inverter_model : inverter_model_record := (multiplier_init_values, init_lcr_model_integrator_gains(5e3, 1000), init_state_variable_gain(500), 0, 0, 0, 0, 0, 4);

------------------------------------------------------------------------
    procedure create_inverter_model (
        signal inverter_model : inout inverter_model_record;
        dc_link_load_current : in int18;
        load_current : in int18);
------------------------------------------------------------------------
    procedure request_inverter_calculation (
        signal inverter_model : out inverter_model_record;
        duty_ratio : in int18);

------------------------------------------------------------------------
end package inverter_model_pkg;

package body inverter_model_pkg is

    procedure create_inverter_model
    (
        signal inverter_model : inout inverter_model_record;
        dc_link_load_current : in int18;
        load_current : in int18
    ) is
        alias inverter_multiplier is inverter_model.inverter_multiplier;
        alias dc_link_voltage is inverter_model.dc_link_voltage;
        alias dc_link_current is inverter_model.dc_link_current;
        alias inverter_lc_filter is inverter_model.inverter_lc_filter;
        alias input_voltage is inverter_model.input_voltage;
        alias grid_inverter_state_counter is inverter_model.grid_inverter_state_counter;
        alias duty_ratio is inverter_model.duty_ratio;

    --------------------------------------------------
        impure function "*" ( left, right : int18)
        return int18
        is
        begin
            sequential_multiply(inverter_multiplier, left, right);
            return get_multiplier_result(inverter_multiplier, 15);
        end "*";
    --------------------------------------------------

    begin
        create_multiplier(inverter_multiplier);
        create_state_variable(dc_link_voltage, inverter_multiplier, -dc_link_current + dc_link_load_current); 
        create_lcr_filter(inverter_lc_filter, inverter_multiplier, input_voltage - inverter_lc_filter.capacitor_voltage, inverter_lc_filter.inductor_current.state - load_current);

        CASE grid_inverter_state_counter is
            WHEN 0 =>
                multiply(inverter_multiplier, dc_link_voltage.state, duty_ratio);
                grid_inverter_state_counter <= grid_inverter_state_counter + 1;
            WHEN 1 =>
                multiply(inverter_multiplier, inverter_lc_filter.inductor_current.state, duty_ratio);
                grid_inverter_state_counter <= grid_inverter_state_counter + 1;
            WHEN 2 =>
                if multiplier_is_ready(inverter_multiplier) then
                    input_voltage <= get_multiplier_result(inverter_multiplier, 15);
                    grid_inverter_state_counter <= grid_inverter_state_counter + 1;
                end if;
            WHEN 3 =>
                dc_link_current <= get_multiplier_result(inverter_multiplier, 15);
                grid_inverter_state_counter <= grid_inverter_state_counter + 1;
            WHEN 4 =>
                calculate(dc_link_voltage);
                increment_counter_when_ready(inverter_multiplier, grid_inverter_state_counter);
            WHEN 5 =>
                calculate_lcr_filter(inverter_lc_filter);
                grid_inverter_state_counter <= grid_inverter_state_counter + 1;
            WHEN others => -- wait for restart
        end CASE;
        
    end create_inverter_model;

------------------------------------------------------------------------
    procedure request_inverter_calculation
    (
        signal inverter_model : out inverter_model_record;
        duty_ratio : in int18
    ) is
    begin
        inverter_model.grid_inverter_state_counter <= 0;
        inverter_model.duty_ratio <= duty_ratio;
    end  request_inverter_calculation;

end package body inverter_model_pkg; 
